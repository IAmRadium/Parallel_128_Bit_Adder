`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:09:50 02/07/2019 
// Design Name: 
// Module Name:    ADD_IMP128_4Bits 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ADD_IMP128_4Bits(a4_1,a4_2,a4_3,a4_4,a4_5,a4_6,a4_7,a4_8,a4_9,a4_10,a4_11,a4_12,a4_13,a4_14,a4_15,a4_16,
a4_17,a4_18,a4_19,a4_20,a4_21,a4_22,a4_23,a4_24,a4_25,a4_26,a4_27,a4_28,a4_29,a4_30,a4_31,a4_32,a4_33,a4_34,a4_35,a4_36,a4_37,a4_38,a4_39,a4_40,
a4_41,a4_42,a4_43,a4_44,a4_45,a4_46,a4_47,a4_48,a4_49,a4_50,a4_51,a4_52,a4_53,a4_54,a4_55,a4_56,a4_57,a4_58,a4_59,a4_60,a4_61,a4_62,a4_63,a4_64,
a4_65,a4_66,a4_67,a4_68,a4_69,a4_70,a4_71,a4_72,a4_73,a4_74,a4_75,a4_76,a4_77,a4_78,a4_79,a4_80,a4_81,a4_82,a4_83,a4_84,a4_85,a4_86,a4_87,a4_88,a4_89,
a4_90,a4_91,a4_92,a4_93,a4_94,a4_95,a4_96,a4_97,a4_98,a4_99,a4_100,a4_101,a4_102,a4_103,a4_104,a4_105,a4_106,a4_107,a4_108,a4_109,a4_110,a4_111,
a4_112,a4_113,a4_114,a4_115,a4_116,a4_117,a4_118,a4_119,a4_120,a4_121,a4_122,a4_123,a4_124,a4_125,a4_126,a4_127,a4_128,
a5_out1,a5_out2,a5_out3,a5_out4,a5_out5,a5_out6,a5_out7,a5_out8,a5_out9,a5_out10,a5_out11,a5_out12,a5_out13,a5_out14,a5_out15,a5_out16,
a5_out17,a5_out18,a5_out19,a5_out20,a5_out21,a5_out22,a5_out23,a5_out24,a5_out25,a5_out26,a5_out27,a5_out28,a5_out29,a5_out30,a5_out31,a5_out32,
a5_out33,a5_out34,a5_out35,a5_out36,a5_out37,a5_out38,a5_out39,a5_out40,a5_out41,a5_out42,a5_out43,a5_out44,a5_out45,a5_out46,a5_out47,a5_out48,
a5_out49,a5_out50,a5_out51,a5_out52,a5_out53,a5_out54,a5_out55,a5_out56,a5_out57,a5_out58,a5_out59,a5_out60,a5_out61,a5_out62,a5_out63,a5_out64);

input [0:3] a4_1,a4_2,a4_3,a4_4,a4_5,a4_6,a4_7,a4_8,a4_9,a4_10,a4_11,a4_12,a4_13,a4_14,a4_15,a4_16,
a4_17,a4_18,a4_19,a4_20,a4_21,a4_22,a4_23,a4_24,a4_25,a4_26,a4_27,a4_28,a4_29,a4_30,a4_31,a4_32,a4_33,a4_34,a4_35,a4_36,a4_37,a4_38,a4_39,a4_40,
a4_41,a4_42,a4_43,a4_44,a4_45,a4_46,a4_47,a4_48,a4_49,a4_50,a4_51,a4_52,a4_53,a4_54,a4_55,a4_56,a4_57,a4_58,a4_59,a4_60,a4_61,a4_62,a4_63,a4_64,
a4_65,a4_66,a4_67,a4_68,a4_69,a4_70,a4_71,a4_72,a4_73,a4_74,a4_75,a4_76,a4_77,a4_78,a4_79,a4_80,a4_81,a4_82,a4_83,a4_84,a4_85,a4_86,a4_87,a4_88,a4_89,
a4_90,a4_91,a4_92,a4_93,a4_94,a4_95,a4_96,a4_97,a4_98,a4_99,a4_100,a4_101,a4_102,a4_103,a4_104,a4_105,a4_106,a4_107,a4_108,a4_109,a4_110,a4_111,
a4_112,a4_113,a4_114,a4_115,a4_116,a4_117,a4_118,a4_119,a4_120,a4_121,a4_122,a4_123,a4_124,a4_125,a4_126,a4_127,a4_128;

output [0:4] a5_out1,a5_out2,a5_out3,a5_out4,a5_out5,a5_out6,a5_out7,a5_out8,a5_out9,a5_out10,a5_out11,a5_out12,a5_out13,a5_out14,a5_out15,a5_out16,
a5_out17,a5_out18,a5_out19,a5_out20,a5_out21,a5_out22,a5_out23,a5_out24,a5_out25,a5_out26,a5_out27,a5_out28,a5_out29,a5_out30,a5_out31,a5_out32,
a5_out33,a5_out34,a5_out35,a5_out36,a5_out37,a5_out38,a5_out39,a5_out40,a5_out41,a5_out42,a5_out43,a5_out44,a5_out45,a5_out46,a5_out47,a5_out48,
a5_out49,a5_out50,a5_out51,a5_out52,a5_out53,a5_out54,a5_out55,a5_out56,a5_out57,a5_out58,a5_out59,a5_out60,a5_out61,a5_out62,a5_out63,a5_out64;


ADD_4Bit a40(.a4(a4_1),.b4(a4_2),.f5(a5_out1));
ADD_4Bit a41(.a4(a4_3),.b4(a4_4),.f5(a5_out2));
ADD_4Bit a42(.a4(a4_5),.b4(a4_6),.f5(a5_out3));
ADD_4Bit a43(.a4(a4_7),.b4(a4_8),.f5(a5_out4));
ADD_4Bit a44(.a4(a4_9),.b4(a4_10),.f5(a5_out5));
ADD_4Bit a45(.a4(a4_11),.b4(a4_12),.f5(a5_out6));
ADD_4Bit a46(.a4(a4_13),.b4(a4_14),.f5(a5_out7));
ADD_4Bit a47(.a4(a4_15),.b4(a4_16),.f5(a5_out8));
ADD_4Bit a48(.a4(a4_17),.b4(a4_18),.f5(a5_out9));
ADD_4Bit a49(.a4(a4_19),.b4(a4_20),.f5(a5_out10));
ADD_4Bit a410(.a4(a4_21),.b4(a4_22),.f5(a5_out11));
ADD_4Bit a411(.a4(a4_23),.b4(a4_24),.f5(a5_out12));
ADD_4Bit a412(.a4(a4_25),.b4(a4_26),.f5(a5_out13));
ADD_4Bit a413(.a4(a4_27),.b4(a4_28),.f5(a5_out14));
ADD_4Bit a414(.a4(a4_29),.b4(a4_30),.f5(a5_out15));
ADD_4Bit a415(.a4(a4_31),.b4(a4_32),.f5(a5_out16));
ADD_4Bit a416(.a4(a4_33),.b4(a4_34),.f5(a5_out17));
ADD_4Bit a417(.a4(a4_35),.b4(a4_36),.f5(a5_out18));
ADD_4Bit a418(.a4(a4_37),.b4(a4_38),.f5(a5_out19));
ADD_4Bit a419(.a4(a4_39),.b4(a4_40),.f5(a5_out20));
ADD_4Bit a420(.a4(a4_41),.b4(a4_42),.f5(a5_out21));
ADD_4Bit a421(.a4(a4_43),.b4(a4_44),.f5(a5_out22));
ADD_4Bit a422(.a4(a4_45),.b4(a4_46),.f5(a5_out23));
ADD_4Bit a423(.a4(a4_47),.b4(a4_48),.f5(a5_out24));
ADD_4Bit a424(.a4(a4_49),.b4(a4_50),.f5(a5_out25));
ADD_4Bit a425(.a4(a4_51),.b4(a4_52),.f5(a5_out26));
ADD_4Bit a426(.a4(a4_53),.b4(a4_54),.f5(a5_out27));
ADD_4Bit a427(.a4(a4_55),.b4(a4_56),.f5(a5_out28));
ADD_4Bit a428(.a4(a4_57),.b4(a4_58),.f5(a5_out29));
ADD_4Bit a429(.a4(a4_59),.b4(a4_60),.f5(a5_out30));
ADD_4Bit a430(.a4(a4_61),.b4(a4_62),.f5(a5_out31));
ADD_4Bit a431(.a4(a4_63),.b4(a4_64),.f5(a5_out32));
ADD_4Bit a432(.a4(a4_65),.b4(a4_66),.f5(a5_out33));
ADD_4Bit a433(.a4(a4_67),.b4(a4_68),.f5(a5_out34));
ADD_4Bit a434(.a4(a4_69),.b4(a4_70),.f5(a5_out35));
ADD_4Bit a435(.a4(a4_71),.b4(a4_72),.f5(a5_out36));
ADD_4Bit a436(.a4(a4_73),.b4(a4_74),.f5(a5_out37));
ADD_4Bit a437(.a4(a4_75),.b4(a4_76),.f5(a5_out38));
ADD_4Bit a438(.a4(a4_77),.b4(a4_78),.f5(a5_out39));
ADD_4Bit a439(.a4(a4_79),.b4(a4_80),.f5(a5_out40));
ADD_4Bit a440(.a4(a4_81),.b4(a4_82),.f5(a5_out41));
ADD_4Bit a441(.a4(a4_83),.b4(a4_84),.f5(a5_out42));
ADD_4Bit a442(.a4(a4_85),.b4(a4_86),.f5(a5_out43));
ADD_4Bit a443(.a4(a4_87),.b4(a4_88),.f5(a5_out44));
ADD_4Bit a444(.a4(a4_89),.b4(a4_90),.f5(a5_out45));
ADD_4Bit a445(.a4(a4_91),.b4(a4_92),.f5(a5_out46));
ADD_4Bit a446(.a4(a4_93),.b4(a4_94),.f5(a5_out47));
ADD_4Bit a447(.a4(a4_95),.b4(a4_96),.f5(a5_out48));
ADD_4Bit a448(.a4(a4_97),.b4(a4_98),.f5(a5_out49));
ADD_4Bit a449(.a4(a4_99),.b4(a4_100),.f5(a5_out50));
ADD_4Bit a450(.a4(a4_101),.b4(a4_102),.f5(a5_out51));
ADD_4Bit a451(.a4(a4_103),.b4(a4_104),.f5(a5_out52));
ADD_4Bit a452(.a4(a4_105),.b4(a4_106),.f5(a5_out53));
ADD_4Bit a453(.a4(a4_107),.b4(a4_108),.f5(a5_out54));
ADD_4Bit a454(.a4(a4_109),.b4(a4_110),.f5(a5_out55));
ADD_4Bit a455(.a4(a4_111),.b4(a4_112),.f5(a5_out56));
ADD_4Bit a456(.a4(a4_113),.b4(a4_114),.f5(a5_out57));
ADD_4Bit a457(.a4(a4_115),.b4(a4_116),.f5(a5_out58));
ADD_4Bit a458(.a4(a4_117),.b4(a4_118),.f5(a5_out59));
ADD_4Bit a459(.a4(a4_119),.b4(a4_120),.f5(a5_out60));
ADD_4Bit a460(.a4(a4_121),.b4(a4_122),.f5(a5_out61));
ADD_4Bit a461(.a4(a4_123),.b4(a4_124),.f5(a5_out62));
ADD_4Bit a462(.a4(a4_125),.b4(a4_126),.f5(a5_out63));
ADD_4Bit a463(.a4(a4_127),.b4(a4_128),.f5(a5_out64));

endmodule
