`timescale 1ns / 1ps
`include "ADD_IMP.v"

module test4_TB;

	// Inputs
	reg [3:0] a1;
	reg [3:0] a2;
	reg [3:0] a3;
	reg [3:0] a4;
	reg [3:0] a5;
	reg [3:0] a6;
	reg [3:0] a7;
	reg [3:0] a8;
	reg [3:0] a9;
	reg [3:0] a10;
	reg [3:0] a11;
	reg [3:0] a12;
	reg [3:0] a13;
	reg [3:0] a14;
	reg [3:0] a15;
	reg [3:0] a16;
	reg [3:0] a17;
	reg [3:0] a18;
	reg [3:0] a19;
	reg [3:0] a20;
	reg [3:0] a21;
	reg [3:0] a22;
	reg [3:0] a23;
	reg [3:0] a24;
	reg [3:0] a25;
	reg [3:0] a26;
	reg [3:0] a27;
	reg [3:0] a28;
	reg [3:0] a29;
	reg [3:0] a30;
	reg [3:0] a31;
	reg [3:0] a32;
	reg [3:0] a33;
	reg [3:0] a34;
	reg [3:0] a35;
	reg [3:0] a36;
	reg [3:0] a37;
	reg [3:0] a38;
	reg [3:0] a39;
	reg [3:0] a40;
	reg [3:0] a41;
	reg [3:0] a42;
	reg [3:0] a43;
	reg [3:0] a44;
	reg [3:0] a45;
	reg [3:0] a46;
	reg [3:0] a47;
	reg [3:0] a48;
	reg [3:0] a49;
	reg [3:0] a50;
	reg [3:0] a51;
	reg [3:0] a52;
	reg [3:0] a53;
	reg [3:0] a54;
	reg [3:0] a55;
	reg [3:0] a56;
	reg [3:0] a57;
	reg [3:0] a58;
	reg [3:0] a59;
	reg [3:0] a60;
	reg [3:0] a61;
	reg [3:0] a62;
	reg [3:0] a63;
	reg [3:0] a64;
	reg [3:0] a65;
	reg [3:0] a66;
	reg [3:0] a67;
	reg [3:0] a68;
	reg [3:0] a69;
	reg [3:0] a70;
	reg [3:0] a71;
	reg [3:0] a72;
	reg [3:0] a73;
	reg [3:0] a74;
	reg [3:0] a75;
	reg [3:0] a76;
	reg [3:0] a77;
	reg [3:0] a78;
	reg [3:0] a79;
	reg [3:0] a80;
	reg [3:0] a81;
	reg [3:0] a82;
	reg [3:0] a83;
	reg [3:0] a84;
	reg [3:0] a85;
	reg [3:0] a86;
	reg [3:0] a87;
	reg [3:0] a88;
	reg [3:0] a89;
	reg [3:0] a90;
	reg [3:0] a91;
	reg [3:0] a92;
	reg [3:0] a93;
	reg [3:0] a94;
	reg [3:0] a95;
	reg [3:0] a96;
	reg [3:0] a97;
	reg [3:0] a98;
	reg [3:0] a99;
	reg [3:0] a100;
	reg [3:0] a101;
	reg [3:0] a102;
	reg [3:0] a103;
	reg [3:0] a104;
	reg [3:0] a105;
	reg [3:0] a106;
	reg [3:0] a107;
	reg [3:0] a108;
	reg [3:0] a109;
	reg [3:0] a110;
	reg [3:0] a111;
	reg [3:0] a112;
	reg [3:0] a113;
	reg [3:0] a114;
	reg [3:0] a115;
	reg [3:0] a116;
	reg [3:0] a117;
	reg [3:0] a118;
	reg [3:0] a119;
	reg [3:0] a120;
	reg [3:0] a121;
	reg [3:0] a122;
	reg [3:0] a123;
	reg [3:0] a124;
	reg [3:0] a125;
	reg [3:0] a126;
	reg [3:0] a127;
	reg [3:0] a128;

	// Outputs
	wire [10:0] a11_out;

	// Instantiate the Unit Under Test (UUT)
	ADD_IMP uut (
		.a1(a1), 
		.a2(a2), 
		.a3(a3), 
		.a4(a4), 
		.a5(a5), 
		.a6(a6), 
		.a7(a7), 
		.a8(a8), 
		.a9(a9), 
		.a10(a10), 
		.a11(a11), 
		.a12(a12), 
		.a13(a13), 
		.a14(a14), 
		.a15(a15), 
		.a16(a16), 
		.a17(a17), 
		.a18(a18), 
		.a19(a19), 
		.a20(a20), 
		.a21(a21), 
		.a22(a22), 
		.a23(a23), 
		.a24(a24), 
		.a25(a25), 
		.a26(a26), 
		.a27(a27), 
		.a28(a28), 
		.a29(a29), 
		.a30(a30), 
		.a31(a31), 
		.a32(a32), 
		.a33(a33), 
		.a34(a34), 
		.a35(a35), 
		.a36(a36), 
		.a37(a37), 
		.a38(a38), 
		.a39(a39), 
		.a40(a40), 
		.a41(a41), 
		.a42(a42), 
		.a43(a43), 
		.a44(a44), 
		.a45(a45), 
		.a46(a46), 
		.a47(a47), 
		.a48(a48), 
		.a49(a49), 
		.a50(a50), 
		.a51(a51), 
		.a52(a52), 
		.a53(a53), 
		.a54(a54), 
		.a55(a55), 
		.a56(a56), 
		.a57(a57), 
		.a58(a58), 
		.a59(a59), 
		.a60(a60), 
		.a61(a61), 
		.a62(a62), 
		.a63(a63), 
		.a64(a64), 
		.a65(a65), 
		.a66(a66), 
		.a67(a67), 
		.a68(a68), 
		.a69(a69), 
		.a70(a70), 
		.a71(a71), 
		.a72(a72), 
		.a73(a73), 
		.a74(a74), 
		.a75(a75), 
		.a76(a76), 
		.a77(a77), 
		.a78(a78), 
		.a79(a79), 
		.a80(a80), 
		.a81(a81), 
		.a82(a82), 
		.a83(a83), 
		.a84(a84), 
		.a85(a85), 
		.a86(a86), 
		.a87(a87), 
		.a88(a88), 
		.a89(a89), 
		.a90(a90), 
		.a91(a91), 
		.a92(a92), 
		.a93(a93), 
		.a94(a94), 
		.a95(a95), 
		.a96(a96), 
		.a97(a97), 
		.a98(a98), 
		.a99(a99), 
		.a100(a100), 
		.a101(a101), 
		.a102(a102), 
		.a103(a103), 
		.a104(a104), 
		.a105(a105), 
		.a106(a106), 
		.a107(a107), 
		.a108(a108), 
		.a109(a109), 
		.a110(a110), 
		.a111(a111), 
		.a112(a112), 
		.a113(a113), 
		.a114(a114), 
		.a115(a115), 
		.a116(a116), 
		.a117(a117), 
		.a118(a118), 
		.a119(a119), 
		.a120(a120), 
		.a121(a121), 
		.a122(a122), 
		.a123(a123), 
		.a124(a124), 
		.a125(a125), 
		.a126(a126), 
		.a127(a127), 
		.a128(a128), 
		.a11_out(a11_out)
	);

	initial begin
		$dumpfile("test4.vcd");
		$dumpvars(0,test4_TB);
		// Initialize Inputs
		a1 = 4'b1111;
		a2 = 4'b1111;
		a3 = 4'b1111;
		a4 = 4'b1111;
		a5 = 4'b1111;
		a6 = 4'b1111;
		a7 = 4'b0001;
		a8 = 4'b0001;
		a9 = 4'b0001;
		a10 = 4'b0001;
		a11 = 4'b0001;
		a12 = 4'b0001;
		a13 = 4'b0001;
		a14 = 4'b0001;
		a15 = 4'b0001;
		a16 = 4'b0001;
		a17 = 4'b0001;
		a18 = 4'b0001;
		a19 = 4'b0001;
		a20 = 4'b0001;
		a21 = 4'b0001;
		a22 = 4'b0001;
		a23 = 4'b0001;
		a24 = 4'b0001;
		a25 = 4'b0001;
		a26 = 4'b0001;
		a27 = 4'b0001;
		a28 = 4'b0001;
		a29 = 4'b0001;
		a30 = 4'b0001;
		a31 = 4'b0001;
		a32 = 4'b0001;
		a33 = 4'b0001;
		a34 = 4'b0001;
		a35 = 4'b0001;
		a36 = 4'b0001;
		a37 = 4'b0001;
		a38 = 4'b0001;
		a39 = 4'b0001;
		a40 = 4'b0001;
		a41 = 4'b0001;
		a42 = 4'b0001;
		a43 = 4'b0001;
		a44 = 4'b0001;
		a45 = 4'b0001;
		a46 = 4'b0001;
		a47 = 4'b0001;
		a48 = 4'b0001;
		a49 = 4'b0001;
		a50 = 4'b0001;
		a51 = 4'b0001;
		a52 = 4'b0001;
		a53 = 4'b0001;
		a54 = 4'b0001;
		a55 = 4'b0001;
		a56 = 4'b0001;
		a57 = 4'b0001;
		a58 = 4'b0001;
		a59 = 4'b0001;
		a60 = 4'b0001;
		a61 = 4'b0001;
		a62 = 4'b0001;
		a63 = 4'b0001;
		a64 = 4'b0001;
		a65 = 4'b0001;
		a66 = 4'b0001;
		a67 = 4'b0001;
		a68 = 4'b0001;
		a69 = 4'b0001;
		a70 = 4'b0001;
		a71 = 4'b0001;
		a72 = 4'b0001;
		a73 = 4'b0001;
		a74 = 4'b0001;
		a75 = 4'b0001;
		a76 = 4'b0001;
		a77 = 4'b0001;
		a78 = 4'b0001;
		a79 = 4'b0001;
		a80 = 4'b0001;
		a81 = 4'b0001;
		a82 = 4'b0001;
		a83 = 4'b0001;
		a84 = 4'b0001;
		a85 = 4'b0001;
		a86 = 4'b0001;
		a87 = 4'b0001;
		a88 = 4'b0001;
		a89 = 4'b0001;
		a90 = 4'b0001;
		a91 = 4'b0001;
		a92 = 4'b0001;
		a93 = 4'b0001;
		a94 = 4'b0001;
		a95 = 4'b0001;
		a96 = 4'b0001;
		a97 = 4'b0001;
		a98 = 4'b0001;
		a99 = 4'b0001;
		a100 = 4'b0001;
		a101 = 4'b0001;
		a102 = 4'b0001;
		a103 = 4'b0001;
		a104 = 4'b0001;
		a105 = 4'b0001;
		a106 = 4'b0001;
		a107 = 4'b0001;
		a108 = 4'b0001;
		a109 = 4'b0001;
		a110 = 4'b0001;
		a111 = 4'b0001;
		a112 = 4'b0001;
		a113 = 4'b0001;
		a114 = 4'b0001;
		a115 = 4'b0001;
		a116 = 4'b0001;
		a117 = 4'b0001;
		a118 = 4'b0001;
		a119 = 4'b0001;
		a120 = 4'b0001;
		a121 = 4'b0001;
		a122 = 4'b0001;
		a123 = 4'b0001;
		a124 = 4'b0001;
		a125 = 4'b0001;
		a126 = 4'b0001;
		a127 = 4'b0001;
		a128 = 4'b0001;


		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

